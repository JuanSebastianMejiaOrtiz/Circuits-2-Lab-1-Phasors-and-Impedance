Lab 1: Phasors and Impedance of the RC Circuit
* Authors: Juan Sebastian Mejia Ortiz, Emmanuel Garces Agudelo

* Voltage Sources
v1 a 0 SIN(0 1 {f} 0 0 90)

* Resistors
r1 a b 1k

* Capacitors
c1 b 0 10nF

* Parameters
.step param f list 2k 20k 200k
.param T = 1/{f}
.param tstart = 0
.param tstop = 2*{T}

* Analysis
.tran 0 {tstop} {tstart}
.end
